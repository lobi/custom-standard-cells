magic
tech sky130A
timestamp 1757244268
<< nwell >>
rect -85 -30 230 65
rect 360 -30 570 65
<< nmos >>
rect 10 -165 35 -110
rect 110 -165 135 -110
rect 440 -165 455 -110
<< pmos >>
rect 10 -10 35 45
rect 110 -10 135 45
rect 440 -10 455 45
<< ndiff >>
rect -65 -135 10 -110
rect -65 -155 -50 -135
rect -30 -155 10 -135
rect -65 -165 10 -155
rect 35 -115 110 -110
rect 35 -135 60 -115
rect 80 -135 110 -115
rect 35 -165 110 -135
rect 135 -135 210 -110
rect 135 -155 175 -135
rect 195 -155 210 -135
rect 135 -165 210 -155
rect 385 -130 440 -110
rect 385 -150 400 -130
rect 420 -150 440 -130
rect 385 -165 440 -150
rect 455 -120 550 -110
rect 455 -140 515 -120
rect 535 -140 550 -120
rect 455 -165 550 -140
<< pdiff >>
rect -65 40 10 45
rect -65 20 -50 40
rect -30 20 10 40
rect -65 -10 10 20
rect 35 -10 110 45
rect 135 20 210 45
rect 135 0 170 20
rect 190 0 210 20
rect 135 -10 210 0
rect 385 30 440 45
rect 385 10 400 30
rect 420 10 440 30
rect 385 -10 440 10
rect 455 25 550 45
rect 455 5 515 25
rect 535 5 550 25
rect 455 -10 550 5
<< ndiffc >>
rect -50 -155 -30 -135
rect 60 -135 80 -115
rect 175 -155 195 -135
rect 400 -150 420 -130
rect 515 -140 535 -120
<< pdiffc >>
rect -50 20 -30 40
rect 170 0 190 20
rect 400 10 420 30
rect 515 5 535 25
<< poly >>
rect 10 45 35 80
rect 110 45 135 80
rect 440 45 455 95
rect 10 -110 35 -10
rect 110 -110 135 -10
rect 287 -45 328 -37
rect 440 -45 455 -10
rect 287 -70 295 -45
rect 320 -70 455 -45
rect 287 -78 328 -70
rect 440 -110 455 -70
rect 10 -185 35 -165
rect 110 -185 135 -165
rect 440 -225 455 -165
<< polycont >>
rect 295 -70 320 -45
<< ndiodelvtc >>
rect 0 95 20 115
rect 105 95 125 115
rect 210 95 230 115
rect 5 -235 25 -215
rect 90 -235 110 -215
rect 200 -235 220 -215
<< locali >>
rect -50 95 0 115
rect 20 95 105 115
rect 125 95 210 115
rect 230 95 420 115
rect -50 40 -30 95
rect -50 5 -30 20
rect 170 20 190 35
rect 170 -45 190 0
rect 400 30 420 95
rect 400 -5 420 10
rect 515 25 535 40
rect 287 -45 328 -37
rect 170 -55 295 -45
rect 60 -70 295 -55
rect 320 -70 328 -45
rect 60 -75 190 -70
rect 60 -115 80 -75
rect 287 -78 328 -70
rect 515 -55 535 5
rect 515 -80 630 -55
rect -50 -135 -30 -125
rect 60 -145 80 -135
rect 175 -135 195 -125
rect -50 -215 -30 -155
rect 175 -215 195 -155
rect 400 -130 420 -115
rect 400 -215 420 -150
rect 515 -120 535 -80
rect 515 -160 535 -140
rect -50 -235 5 -215
rect 25 -235 90 -215
rect 110 -235 200 -215
rect 220 -235 420 -215
<< labels >>
rlabel locali -15 100 -15 100 1 VDD
port 4 n
rlabel locali -25 -225 -25 -225 1 GND
port 3 n
rlabel poly 20 -50 20 -50 1 A
port 1 n
rlabel poly 120 -50 120 -50 1 B
port 2 n
rlabel locali 630 -65 630 -65 7 Y
port 5 w
<< end >>
