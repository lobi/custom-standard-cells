magic
tech sky130A
timestamp 1752848002
<< nwell >>
rect -110 90 300 235
<< nmos >>
rect 10 -50 25 55
rect 215 -50 230 55
<< pmos >>
rect 10 110 25 215
rect 215 110 230 215
<< ndiff >>
rect -40 40 10 55
rect -40 -35 -25 40
rect -5 -35 10 40
rect -40 -50 10 -35
rect 25 40 75 55
rect 25 -35 40 40
rect 60 -35 75 40
rect 25 -50 75 -35
rect 165 40 215 55
rect 165 -35 180 40
rect 200 -35 215 40
rect 165 -50 215 -35
rect 230 40 280 55
rect 230 -35 245 40
rect 265 -35 280 40
rect 230 -50 280 -35
<< pdiff >>
rect -40 200 10 215
rect -40 125 -25 200
rect -5 125 10 200
rect -40 110 10 125
rect 25 200 75 215
rect 25 125 40 200
rect 60 125 75 200
rect 25 110 75 125
rect 165 200 215 215
rect 165 125 180 200
rect 200 125 215 200
rect 165 110 215 125
rect 230 200 280 215
rect 230 125 245 200
rect 265 125 280 200
rect 230 110 280 125
<< ndiffc >>
rect -25 -35 -5 40
rect 40 -35 60 40
rect 180 -35 200 40
rect 245 -35 265 40
<< pdiffc >>
rect -25 125 -5 200
rect 40 125 60 200
rect 180 125 200 200
rect 245 125 265 200
<< psubdiff >>
rect -90 40 -40 55
rect -90 -35 -75 40
rect -55 -35 -40 40
rect -90 -50 -40 -35
rect 115 40 165 55
rect 115 -35 130 40
rect 150 -35 165 40
rect 115 -50 165 -35
<< nsubdiff >>
rect -90 200 -40 215
rect -90 125 -75 200
rect -55 125 -40 200
rect -90 110 -40 125
rect 115 200 165 215
rect 115 125 130 200
rect 150 125 165 200
rect 115 110 165 125
<< psubdiffcont >>
rect -75 -35 -55 40
rect 130 -35 150 40
<< nsubdiffcont >>
rect -75 125 -55 200
rect 130 125 150 200
<< poly >>
rect 10 215 25 230
rect 215 215 230 230
rect 10 55 25 110
rect 215 55 230 110
rect 10 -65 25 -50
rect 215 -65 230 -50
rect -15 -75 25 -65
rect -15 -95 -5 -75
rect 15 -95 25 -75
rect -15 -105 25 -95
rect 190 -75 230 -65
rect 190 -95 200 -75
rect 220 -95 230 -75
rect 190 -105 230 -95
<< polycont >>
rect -5 -95 15 -75
rect 200 -95 220 -75
<< locali >>
rect -85 200 5 210
rect -85 125 -75 200
rect -55 125 -25 200
rect -5 125 5 200
rect -85 115 5 125
rect 30 200 70 210
rect 30 125 40 200
rect 60 125 70 200
rect 30 115 70 125
rect 120 200 210 210
rect 120 125 130 200
rect 150 125 180 200
rect 200 125 210 200
rect 120 115 210 125
rect 235 200 275 210
rect 235 125 245 200
rect 265 125 275 200
rect 235 115 275 125
rect 50 50 70 115
rect 255 50 275 115
rect -85 40 5 50
rect -85 -35 -75 40
rect -55 -35 -25 40
rect -5 -35 5 40
rect -85 -45 5 -35
rect 30 40 70 50
rect 30 -35 40 40
rect 60 -35 70 40
rect 30 -45 70 -35
rect 120 40 210 50
rect 120 -35 130 40
rect 150 -35 180 40
rect 200 -35 210 40
rect 120 -45 210 -35
rect 235 40 275 50
rect 235 -35 245 40
rect 265 -35 275 40
rect 235 -45 275 -35
rect 50 -65 70 -45
rect 255 -65 275 -45
rect -110 -75 25 -65
rect -110 -85 -5 -75
rect -15 -95 -5 -85
rect 15 -95 25 -75
rect 50 -75 230 -65
rect 50 -85 200 -75
rect -15 -105 25 -95
rect 190 -95 200 -85
rect 220 -95 230 -75
rect 255 -85 300 -65
rect 190 -105 230 -95
<< viali >>
rect -75 125 -55 200
rect -25 125 -5 200
rect 130 125 150 200
rect 180 125 200 200
rect -75 -35 -55 40
rect -25 -35 -5 40
rect 130 -35 150 40
rect 180 -35 200 40
<< metal1 >>
rect -110 200 300 210
rect -110 125 -75 200
rect -55 125 -25 200
rect -5 125 130 200
rect 150 125 180 200
rect 200 125 300 200
rect -110 115 300 125
rect -110 40 300 50
rect -110 -35 -75 40
rect -55 -35 -25 40
rect -5 -35 130 40
rect 150 -35 180 40
rect 200 -35 300 40
rect -110 -45 300 -35
<< labels >>
rlabel locali -110 -75 -110 -75 7 A
port 1 w
rlabel metal1 -110 163 -110 163 7 VP
port 3 w
rlabel metal1 -110 2 -110 2 7 VN
port 4 w
rlabel locali 300 -75 300 -75 7 Y
port 2 w
<< end >>
