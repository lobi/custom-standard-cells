magic
tech sky130A
timestamp 1757238157
<< nwell >>
rect -85 0 265 105
<< nmos >>
rect 10 -165 35 -110
rect 145 -165 170 -110
<< pmos >>
rect 10 20 35 75
rect 145 20 170 75
<< ndiff >>
rect -65 -135 10 -110
rect -65 -155 -50 -135
rect -30 -155 10 -135
rect -65 -165 10 -155
rect 35 -125 145 -110
rect 35 -145 60 -125
rect 80 -145 145 -125
rect 35 -165 145 -145
rect 170 -115 245 -110
rect 170 -135 200 -115
rect 220 -135 245 -115
rect 170 -165 245 -135
<< pdiff >>
rect -65 70 10 75
rect -65 50 -50 70
rect -30 50 10 70
rect -65 20 10 50
rect 35 50 145 75
rect 35 30 60 50
rect 80 30 145 50
rect 35 20 145 30
rect 170 70 245 75
rect 170 50 195 70
rect 215 50 245 70
rect 170 20 245 50
<< ndiffc >>
rect -50 -155 -30 -135
rect 60 -145 80 -125
rect 200 -135 220 -115
<< pdiffc >>
rect -50 50 -30 70
rect 60 30 80 50
rect 195 50 215 70
<< poly >>
rect 10 75 35 95
rect 145 75 170 95
rect 10 -35 35 20
rect 145 -10 170 20
rect -30 -45 35 -35
rect -30 -65 -20 -45
rect 0 -65 35 -45
rect 105 -20 170 -10
rect 105 -40 115 -20
rect 135 -40 170 -20
rect 105 -50 170 -40
rect -30 -75 35 -65
rect 10 -110 35 -75
rect 145 -110 170 -50
rect 10 -185 35 -165
rect 145 -185 170 -165
<< polycont >>
rect -20 -65 0 -45
rect 115 -40 135 -20
<< ndiodelvtc >>
rect -65 110 -45 130
rect 0 110 20 130
rect 75 110 95 130
rect 165 110 185 130
rect 225 110 245 130
rect -50 -220 -30 -200
rect 5 -220 25 -200
rect 75 -220 95 -200
rect 165 -220 185 -200
rect 220 -220 240 -200
<< locali >>
rect -85 110 -65 130
rect -45 110 0 130
rect 20 110 75 130
rect 95 110 165 130
rect 185 110 225 130
rect 245 110 265 130
rect -85 105 265 110
rect -50 70 -30 105
rect 195 70 215 105
rect -50 35 -30 50
rect 60 50 80 65
rect 195 35 215 50
rect -30 -45 10 -35
rect -30 -65 -20 -45
rect 0 -65 10 -45
rect -30 -75 10 -65
rect 60 -70 80 30
rect 105 -20 145 -10
rect 105 -40 115 -20
rect 135 -40 145 -20
rect 105 -50 145 -40
rect 60 -90 265 -70
rect 60 -125 80 -90
rect -50 -135 -30 -125
rect 200 -115 220 -90
rect 200 -145 220 -135
rect 60 -155 80 -145
rect -50 -195 -30 -155
rect -85 -200 265 -195
rect -85 -220 -50 -200
rect -30 -220 5 -200
rect 25 -220 75 -200
rect 95 -220 165 -200
rect 185 -220 220 -200
rect 240 -220 265 -200
<< labels >>
rlabel poly 20 -50 20 -50 1 A
port 1 n
rlabel locali -15 115 -15 115 1 VDD
port 5 n
rlabel poly 155 -50 155 -50 1 B
port 2 n
rlabel locali -25 -210 -25 -210 1 GND
port 4 n
rlabel locali 265 -80 265 -80 7 Y
port 3 w
<< end >>
